module module0(
  input   m_clock,
  input   p_reset
);
endmodule
