module module1(
  input   m_clock,
  input   p_reset,
  input   in,
  output  out
);
  assign out = in;
endmodule
