module module0(
  input   in
);
endmodule
