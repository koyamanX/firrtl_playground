module module1(
  input   in,
  output  out
);
  assign out = in;
endmodule
